`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Com
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module orgate(
    input logic a,
    input logic b,
    output logic f

    );
    
    //OR gate
    and u_or(f,a,b);
    
endmodule
